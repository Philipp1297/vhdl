LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY halfadder_test IS
END halfadder_test;

